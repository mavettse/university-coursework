module binario_bcd(bin, dezena, unidade);
	input [4:0] bin;
	output [3:0] dezena, unidade;