module TOPsomador4bits(SW, HEX0, HEX1);
	input [17:0] SW;
	output [6:0] HEX0, HEX1;
		
	wire [3:0] A, B;
	wire TE0;
	
	assign A = SW[17:14];
	assign B = SW[3:0];
	assign TE0 = SW[9];
	
	wire [4:0] S;
	wire [3:0] bcd_unidade, bcd_dezena;
	
	// somador4bits  (a, b, te0,  s);
	somador4bits soma(A, B, TE0, S);

	
	
endmodule